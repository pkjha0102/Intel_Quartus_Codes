module and_gate(out, a, b);
output out;
input a, b;
assign out = a&b;
endmodule

